module tb;
  reg [10:0] a;
  reg [10:0]b;

  initial begin
    $dumpfile("waveform.vcd"); // For GTKWave
    $dumpvars(0, tb);
     a = 11'b00000000000; #10;
     b = 11'b00000000000; #10;
    
    
    // Test pattern 1
    //H                  //H 
    a = 11'b00000000000; b=11'b00000000000;#10;
    a = 11'b11111111111; b=11'b11111111111;#10;
    a = 11'b00000100000; b=11'b00000100000;#10;
    a = 11'b00000100000; b=11'b00000100000;#10;
    a = 11'b00000100000; b=11'b00000100000;#10;
    a = 11'b11111111111; b=11'b11111111111;#10;
    a = 11'b00000000000; b=11'b00000000000;#10;

    // Test pattern 2
    //A                  //E
    a = 11'b00000000000; b= 11'b00000000000;#10;
    a = 11'b00111111111; b= 11'b11111111111;#10;
    a = 11'b01000100000; b= 11'b10000100001;#10;
    a = 11'b10000100000; b= 11'b10000100001;#10;
    a = 11'b01000100000; b= 11'b10000100001;#10;
    a = 11'b00111111111; b= 11'b10000100001;#10;
    a = 11'b00000000000; b= 11'b00000000000;#10;
    
    //R                  //M
    a = 11'b00000000000; b=11'b00000000000; #10;
    a = 11'b11111111111; b=11'b11111111111;#10;
    a = 11'b10000011000; b=11'b01000000000;#10;
    a = 11'b10000010100; b=11'b0110000000;#10;
    a = 11'b10000010010; b=11'b01000000000;#10;
    a = 11'b01111110001; b=11'b11111111111;#10;  // ✅ FIXED: Missing semicolon added
    a = 11'b00000000000; b=11'b00000000000;#10;
    
    //I                   //A
    // Test pattern 3 (Box with center bar)
    a = 11'b00000000000;  b = 11'b00000000000;#10;
    a = 11'b10000000001;  b = 11'b00111111111;#10;
    a = 11'b10000000001;  b = 11'b01000100000;#10;
    a = 11'b10000000001;  b = 11'b10000100000;#10;
    a = 11'b11111111111;  b = 11'b01000100000;#10;
    a = 11'b10000000001;  b = 11'b00100100000;#10;
    a = 11'b10000000001;  b = 11'b00011111111;#10;
    a = 11'b00000000000;  b = 11'b00000000000;#10;
    //N
    b=11'b00000000000;#10;
    b=11'b11111111111;#10;
    b=11'b00111000000;#10;
    b=11'b00000111000;#10;
    b=11'b00000000110;#10;
    b=11'b11111111111;#10;
    b=11'b00000000000;#10;
    
    //T
    b=11'b00000000000;#10;
    b=11'b10000000000;#10;
    b=11'b10000000000;#10;
    b=11'b11111111111;#10;
    b=11'b10000000000;#10;
    b=11'b10000000000;#10;
    b=11'b00000000000;#10;
    
    //H
    b=11'b0000_0000_000;#10;
    b=11'b1111_1111_111;#10;
    b=11'b00000100000;#10;
    b=11'b00000100000;#10;
    b=11'b00000100000;#10;
    b=11'b1111_1111_111;#10;
    b=11'b0000_0000_000;#10;

    $finish;
  end
endmodule
