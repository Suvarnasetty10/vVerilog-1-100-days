//SUVARNA//
module tb;
  reg [10:0]a;
  initial begin
  
    a=11'b00000000000;#10;
    a=11'b11111100001;#10;
    a=11'b10000100001;#10;
    a=11'b10000100001;#10;//Letter S
    a=11'b10000100001;#10;
    a=11'b10000111111;#10;
    a=11'b0000_0000_000;#10;
 
  
    a=11'b00000000000;#10;
    a=11'b11111111111;#10;
    a=11'b00000000001;#10;
    a=11'b00000000001;#10;//letter U
    a=11'b00000000001;#10;
    a=11'b11111111111;#10;
    a=11'b0000_0000_000;#10;
    
    
    a=11'b00000000000;#10;
    a=11'b11111111100;#10;
    a=11'b00000000010;#10;
    a=11'b00000000001;#10;//letter V
    a=11'b00000000010;#10;
    a=11'b11111111100;#10;
    a=11'b0000_0000_000;#10;


    
    a = 11'b00000000000; #10;
    a = 11'b00111111111; #10;
    a = 11'b01000100000; #10;
    a = 11'b10000100000; #10;//letter A
    a = 11'b01000100000; #10;
    a = 11'b00111111111; #10;
    a = 11'b00000000000; #10;
    
    a = 11'b00000000000; #10;
    a = 11'b11111111111;#10;
    a = 11'b10000011000;#10;//letter R
    a = 11'b10000010100;#10;
    a = 11'b10000010010;#10;
    a = 11'b01111110001;#10;  
    a = 11'b00000000000;#10
    
    a=11'b00000000000;#10;
    a=11'b11111111111;#10;
    a=11'b00111000000;#10;
    a=11'b00000111000;#10;//letter N
    a=11'b00000000110;#10;
    a=11'b11111111111;#10;
    a=11'b00000000000;#10;
    
    a = 11'b00000000000; #10;
    a = 11'b00111111111; #10;
    a = 11'b01000100000; #10;
    a = 11'b10000100000; #10;//leeter A
    a = 11'b01000100000; #10;
    a = 11'b00111111111; #10;
    a = 11'b00000000000; #10;
    
  
    
    $finish;
  end
endmodule
